/////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////
`timescale 1ns/1ps
module tb_design();
	
////////////////////////////////////////////////////////////
//参数定义

`define CLK_PERIORD		10		//时钟周期设置为10ns（100MHz）	

////////////////////////////////////////////////////////////
//接口申明

reg a,b,c,d;
reg s0,s1;
wire y;

////////////////////////////////////////////////////////////	
//对被测试的设计进行例化
	
ex1  uut(
        .a(a),
        .b(b),
        .c(c),
        .d(d),
        .s0(s0),
        .s1(s1),
        .y(y)
    );	
	

////////////////////////////////////////////////////////////
//测试激励产生

initial begin
    {a,b,c,d,s0,s1} = 6'b100000;
    #100;
    {a,b,c,d,s0,s1} = 6'b100001;
    #100;
    {a,b,c,d,s0,s1} = 6'b100010;
    #100;
    {a,b,c,d,s0,s1} = 6'b100011;
    #100;

    {a,b,c,d,s0,s1} = 6'b010000;
    #100;
    {a,b,c,d,s0,s1} = 6'b010001;
    #100;
    {a,b,c,d,s0,s1} = 6'b010010;
    #100;
    {a,b,c,d,s0,s1} = 6'b010011;
    #100;

    {a,b,c,d,s0,s1} = 6'b001000;
    #100;
    {a,b,c,d,s0,s1} = 6'b001001;
    #100;
    {a,b,c,d,s0,s1} = 6'b001010;
    #100;
    {a,b,c,d,s0,s1} = 6'b001011;
    #100;

    {a,b,c,d,s0,s1} = 6'b000100;
    #100;
    {a,b,c,d,s0,s1} = 6'b000101;
    #100;
    {a,b,c,d,s0,s1} = 6'b000110;
    #100;
    {a,b,c,d,s0,s1} = 6'b000111;
    #100;

	$stop;
end


endmodule






